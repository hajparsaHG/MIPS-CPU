/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : mul_func                                                     **
 **                                                                          **
 *****************************************************************************/

module mul_func( a,
                 b,
                 clk,
                 hi,
                 lo );

   /*******************************************************************************
   ** The inputs are defined here                                                **
   *******************************************************************************/
   input [31:0] a;
   input [31:0] b;
   input        clk;

   /*******************************************************************************
   ** The outputs are defined here                                               **
   *******************************************************************************/
   output [31:0] hi;
   output [31:0] lo;

   /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
   wire [31:0] s_logisimBus0;
   wire [31:0] s_logisimBus1;
   wire [31:0] s_logisimBus2;
   wire [31:0] s_logisimBus3;

   /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

   /*******************************************************************************
   ** Here all input connections are defined                                     **
   *******************************************************************************/
   assign s_logisimBus0[31:0] = a;
   assign s_logisimBus2[31:0] = b;

   /*******************************************************************************
   ** Here all output connections are defined                                    **
   *******************************************************************************/
   assign hi = s_logisimBus3[31:0];
   assign lo = s_logisimBus1[31:0];

   /*******************************************************************************
   ** Here all normal components are defined                                     **
   *******************************************************************************/
   Multiplier #(.calcBits(64),
                .nrOfBits(32),
                .unsignedMultiplier(0))
      ARITH_1 (.carryIn(32'd0),
               .inputA(s_logisimBus0[31:0]),
               .inputB(s_logisimBus2[31:0]),
               .multHigh(s_logisimBus3[31:0]),
               .multLow(s_logisimBus1[31:0]));


endmodule
